library IEEE;
use IEEE.numeric_std.all;
use IEEE.std_logic_1164.all;

package display_comp is
    constant TEXT_WIDTH      : natural := 80;
    constant TEXT_HEIGHT     : natural := 60;
    constant TILE_WIDTH      : natural := 8;
    constant TILE_HEIGHT     : natural := 8;
    constant PRINTABLE_START : natural := 32;
    constant PRINTABLE_END   : natural := 127;
    constant PRINTABLE_COUNT : natural := PRINTABLE_END - PRINTABLE_START + 1;

    function printable(index : natural) return natural;

    subtype character_t is natural range PRINTABLE_START to PRINTABLE_END;
    type    line_t      is array (0 to TEXT_WIDTH  - 1) of character_t;
    type    glyph_t     is array (0 to 7)               of std_logic_vector(7 downto 0);
    type    glyph_rom_t is array (0 to 127)             of glyph_t;

    constant FONT_ROM : glyph_rom_t := (
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00011000","00111100","00111100","00011000","00011000","00000000","00011000","00000000"),
        ("01101100","01101100","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("01101100","01101100","11111110","01101100","11111110","01101100","01101100","00000000"),
        ("00110000","01111100","11000000","01111000","00001100","11111000","00110000","00000000"),
        ("00000000","11000110","11001100","00011000","00110000","01100110","11000110","00000000"),
        ("00111000","01101100","00111000","01110110","11011100","11001100","01110110","00000000"),
        ("01100000","01100000","11000000","00000000","00000000","00000000","00000000","00000000"),
        ("00011000","00110000","01100000","01100000","01100000","00110000","00011000","00000000"),
        ("01100000","00110000","00011000","00011000","00011000","00110000","01100000","00000000"),
        ("00000000","01100110","00111100","11111111","00111100","01100110","00000000","00000000"),
        ("00000000","00110000","00110000","11111100","00110000","00110000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00110000","00110000","01100000"),
        ("00000000","00000000","00000000","11111100","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00110000","00110000","00000000"),
        ("00000110","00001100","00011000","00110000","01100000","11000000","10000000","00000000"),
        ("01111100","11000110","11001110","11011110","11110110","11100110","01111100","00000000"),
        ("00110000","01110000","00110000","00110000","00110000","00110000","11111100","00000000"),
        ("01111000","11001100","00001100","00111000","01100000","11001100","11111100","00000000"),
        ("01111000","11001100","00001100","00111000","00001100","11001100","01111000","00000000"),
        ("00011100","00111100","01101100","11001100","11111110","00001100","00011110","00000000"),
        ("11111100","11000000","11111000","00001100","00001100","11001100","01111000","00000000"),
        ("00111000","01100000","11000000","11111000","11001100","11001100","01111000","00000000"),
        ("11111100","11001100","00001100","00011000","00110000","00110000","00110000","00000000"),
        ("01111000","11001100","11001100","01111000","11001100","11001100","01111000","00000000"),
        ("01111000","11001100","11001100","01111100","00001100","00011000","01110000","00000000"),
        ("00000000","00110000","00110000","00000000","00000000","00110000","00110000","00000000"),
        ("00000000","00110000","00110000","00000000","00000000","00110000","00110000","01100000"),
        ("00011000","00110000","01100000","11000000","01100000","00110000","00011000","00000000"),
        ("00000000","00000000","11111100","00000000","00000000","11111100","00000000","00000000"),
        ("01100000","00110000","00011000","00001100","00011000","00110000","01100000","00000000"),
        ("01111000","11001100","00001100","00011000","00110000","00000000","00110000","00000000"),
        ("01111100","11000110","11011110","11011110","11011110","11000000","01111000","00000000"),
        ("00110000","01111000","11001100","11001100","11111100","11001100","11001100","00000000"),
        ("11111100","01100110","01100110","01111100","01100110","01100110","11111100","00000000"),
        ("00111100","01100110","11000000","11000000","11000000","01100110","00111100","00000000"),
        ("11111000","01101100","01100110","01100110","01100110","01101100","11111000","00000000"),
        ("11111110","01100010","01101000","01111000","01101000","01100010","11111110","00000000"),
        ("11111110","01100010","01101000","01111000","01101000","01100000","11110000","00000000"),
        ("00111100","01100110","11000000","11000000","11001110","01100110","00111110","00000000"),
        ("11001100","11001100","11001100","11111100","11001100","11001100","11001100","00000000"),
        ("01111000","00110000","00110000","00110000","00110000","00110000","01111000","00000000"),
        ("00011110","00001100","00001100","00001100","11001100","11001100","01111000","00000000"),
        ("11100110","01100110","01101100","01111000","01101100","01100110","11100110","00000000"),
        ("11110000","01100000","01100000","01100000","01100010","01100110","11111110","00000000"),
        ("11000110","11101110","11111110","11111110","11010110","11000110","11000110","00000000"),
        ("11000110","11100110","11110110","11011110","11001110","11000110","11000110","00000000"),
        ("00111000","01101100","11000110","11000110","11000110","01101100","00111000","00000000"),
        ("11111100","01100110","01100110","01111100","01100000","01100000","11110000","00000000"),
        ("01111000","11001100","11001100","11001100","11011100","01111000","00011100","00000000"),
        ("11111100","01100110","01100110","01111100","01101100","01100110","11100110","00000000"),
        ("01111000","11001100","11100000","01110000","00011100","11001100","01111000","00000000"),
        ("11111100","10110100","00110000","00110000","00110000","00110000","01111000","00000000"),
        ("11001100","11001100","11001100","11001100","11001100","11001100","11111100","00000000"),
        ("11001100","11001100","11001100","11001100","11001100","01111000","00110000","00000000"),
        ("11000110","11000110","11000110","11010110","11111110","11101110","11000110","00000000"),
        ("11000110","11000110","01101100","00111000","00111000","01101100","11000110","00000000"),
        ("11001100","11001100","11001100","01111000","00110000","00110000","01111000","00000000"),
        ("11111110","11000110","10001100","00011000","00110010","01100110","11111110","00000000"),
        ("01111000","01100000","01100000","01100000","01100000","01100000","01111000","00000000"),
        ("11000000","01100000","00110000","00011000","00001100","00000110","00000010","00000000"),
        ("01111000","00011000","00011000","00011000","00011000","00011000","01111000","00000000"),
        ("00010000","00111000","01101100","11000110","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111111"),
        ("00110000","00110000","00011000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","01111000","00001100","01111100","11001100","01110110","00000000"),
        ("11100000","01100000","01100000","01111100","01100110","01100110","11011100","00000000"),
        ("00000000","00000000","01111000","11001100","11000000","11001100","01111000","00000000"),
        ("00011100","00001100","00001100","01111100","11001100","11001100","01110110","00000000"),
        ("00000000","00000000","01111000","11001100","11111100","11000000","01111000","00000000"),
        ("00111000","01101100","01100000","11110000","01100000","01100000","11110000","00000000"),
        ("00000000","00000000","01110110","11001100","11001100","01111100","00001100","11111000"),
        ("11100000","01100000","01101100","01110110","01100110","01100110","11100110","00000000"),
        ("00110000","00000000","01110000","00110000","00110000","00110000","01111000","00000000"),
        ("00001100","00000000","00001100","00001100","00001100","11001100","11001100","01111000"),
        ("11100000","01100000","01100110","01101100","01111000","01101100","11100110","00000000"),
        ("01110000","00110000","00110000","00110000","00110000","00110000","01111000","00000000"),
        ("00000000","00000000","11001100","11111110","11111110","11010110","11000110","00000000"),
        ("00000000","00000000","11111000","11001100","11001100","11001100","11001100","00000000"),
        ("00000000","00000000","01111000","11001100","11001100","11001100","01111000","00000000"),
        ("00000000","00000000","11011100","01100110","01100110","01111100","01100000","11110000"),
        ("00000000","00000000","01110110","11001100","11001100","01111100","00001100","00011110"),
        ("00000000","00000000","11011100","01110110","01100110","01100000","11110000","00000000"),
        ("00000000","00000000","01111100","11000000","01111000","00001100","11111000","00000000"),
        ("00010000","00110000","01111100","00110000","00110000","00110100","00011000","00000000"),
        ("00000000","00000000","11001100","11001100","11001100","11001100","01110110","00000000"),
        ("00000000","00000000","11001100","11001100","11001100","01111000","00110000","00000000"),
        ("00000000","00000000","11000110","11010110","11111110","11111110","01101100","00000000"),
        ("00000000","00000000","11000110","01101100","00111000","01101100","11000110","00000000"),
        ("00000000","00000000","11001100","11001100","11001100","01111100","00001100","11111000"),
        ("00000000","00000000","11111100","10011000","00110000","01100100","11111100","00000000"),
        ("00011100","00110000","00110000","11100000","00110000","00110000","00011100","00000000"),
        ("00011000","00011000","00011000","00000000","00011000","00011000","00011000","00000000"),
        ("11100000","00110000","00110000","00011100","00110000","00110000","11100000","00000000"),
        ("01110110","11011100","00000000","00000000","00000000","00000000","00000000","00000000"),
        ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"));

end package;

package body display_comp is
    function printable(index : natural) return natural is
    begin
        return PRINTABLE_START + index;
    end function;
end package body;
